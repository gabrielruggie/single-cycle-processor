module MemoryWriteBackRegister ();



endmodule