module WriteBackStage ();

    // 1. Choose between ALU or Memory output to write back
        // Remember enable on the register file will dictate if this matters

endmodule