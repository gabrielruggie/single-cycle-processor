module DecodeExecuteRegister (

    

);




endmodule