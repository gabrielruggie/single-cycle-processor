module ExecuteStage ();

    // 1. ALU Input Logic
    
    // 2. Register Value Logic

    // 3. ALU

    // 4. Data Hazard Unit

endmodule