module DecodeStage ();

    // 1. Register File

    // 2. Control Unit

    // 3. Flag Register

    // 4. Control Hazard Unit

    // 5. Register & Imm. Dataflow

    // 6. Stalls & Flush Logic

endmodule