module FetchStage ();

    // 1. Calculate PC Halt

    // 2. PC Control Unit In

    // 3. PC Register

    // 4. Instruction Memory

    // 5. PC Control Unit

endmodule