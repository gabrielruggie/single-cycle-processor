module MemoryStage ();

    // 1. Logic to determine inputs

    // 2. Data Memory
    
endmodule