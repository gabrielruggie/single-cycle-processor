module ControlHazardUnit (



);

endmodule