module ExecuteMemoryRegister ();



endmodule