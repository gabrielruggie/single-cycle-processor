module (

    input [3:0] opcode,
    output dst_reg, alu_src, mem_read, mem_write, mem_to_reg, write_reg, branch_en, branch, pcs, lower_half, upper_half;

);

    reg _dst_reg, _alu_src, _mem_read, _mem_write, _mem_to_reg, _write_reg, _branch_en, _branch, _pcs, _lower_half, _upper_half;

    assign 

endmodule