module DataHazardUnit (

    

);

endmodule